PrimarySMTPAddress
jmarton@hsc.wvu.edu
pmartone@hsc.wvu.edu
mamonahan-Retired@hsc.wvu.edu
mzeppuhar-retiree@WVUHSC.onmicrosoft.com
nancy.marzella@hsc.wvu.edu
tamashburn@hsc.wvu.edu
acmason@hsc.wvu.edu
jdmason@hsc.wvu.edu
kmason@hsc.wvu.edu
michael.mason@hsc.wvu.edu
jmassie@hsc.wvu.edu
AMASSOUD@hsc.wvu.edu
fmastalerz@hsc.wvu.edu
fmatalkah@hsc.wvu.edu
KMMATHAI@hsc.wvu.edu
adriane.matheny@hsc.wvu.edu
hmatheny@hsc.wvu.edu
pmathers@hsc.wvu.edu
pmathew@WVUHSC.onmicrosoft.com
rmathews@hsc.wvu.edu
tmatlick@hsc.wvu.edu
JAMATONAK@hsc.wvu.edu
mamatos@hsc.wvu.edu
mamattagonzalez@hsc.wvu.edu
rsmatteotti@hsc.wvu.edu
mdmattes@hsc.wvu.edu
chelsi.matthews@hsc.wvu.edu
jknox3@hsc.wvu.edu
matthewsjproxywvuh@WVUHSC.onmicrosoft.com
Amy.Matuga@hsc.wvu.edu
irene.maundu@hsc.wvu.edu
KDMAUPIN@hsc.wvu.edu
MAMAURER@hsc.wvu.edu
mmawhinney@hsc.wvu.edu
crmay@hsc.wvu.edu
mmayfield@hsc.wvu.edu
tmayfield@hsc.wvu.edu
Chasity.Mayhew@hsc.wvu.edu
camayhew@hsc.wvu.edu
jamayle@hsc.wvu.edu
lmayle@hsc.wvu.edu
slmayle@hsc.wvu.edu
chmaynard@hsc.wvu.edu
lmaynor@hsc.wvu.edu
rmayolo@hsc.wvu.edu
khurt@hsc.wvu.edu
dmazon1@hsc.wvu.edu
jmazza@hsc.wvu.edu
bjm0039@hsc.wvu.edu
gmmazzetti@hsc.wvu.edu
MBRCC_1612@hsc.wvu.edu
rmcgahan@hsc.wvu.edu
jmmcbee@hsc.wvu.edu
kimberly.mcbrayer@hsc.wvu.edu
cmcbride@hsc.wvu.edu
cmcburney@hsc.wvu.edu
mccabebproxywvuh@WVUHSC.onmicrosoft.com
jamie.mccall@hsc.wvu.edu
KYMCCALLISTER@hsc.wvu.edu
tdmccallister@hsc.wvu.edu
kmccammon@hsc.wvu.edu
lmccartney@hsc.wvu.edu
dmccarty@hsc.wvu.edu
mamccawley@hsc.wvu.edu
jmcchesney@hsc.wvu.edu
rmcclai4@hsc.wvu.edu
djmcclelland@hsc.wvu.edu
ryan.mccloy@hsc.wvu.edu
kevin.mccluskey@hsc.wvu.edu
rmccluskey@hsc.wvu.edu
rmccombie@hsc.wvu.edu
bmccormick@hsc.wvu.edu
kamccormick@hsc.wvu.edu
william.mccormick1@hsc.wvu.edu
kmccourt@hsc.wvu.edu
tmccourt@hsc.wvu.edu
gmccoy@hsc.wvu.edu
ashley.mccracken@hsc.wvu.edu
amhuckins@hsc.wvu.edu
smccrone@hsc.wvu.edu
jlmccrory@hsc.wvu.edu
cmccross@hsc.wvu.edu
megan.mccullough@hsc.wvu.edu
llmccune@hsc.wvu.edu
pmcdade@hsc.wvu.edu
david.mcdermott@hsc.wvu.edu
PWMCDEVITT@hsc.wvu.edu
mmcdilda@hsc.wvu.edu
bmlong@hsc.wvu.edu
rmcdonald@hsc.wvu.edu
dmcdonnell@hsc.wvu.edu
bmcdonough@hsc.wvu.edu
megan.mcdougal@hsc.wvu.edu
bmcelfis@hsc.wvu.edu
michele.mcelroy@hsc.wvu.edu
smcewuen@hsc.wvu.edu
anthony.mcfarlane@wvumedicine.org
lem00280747@WVUHSC.onmicrosoft.com
dmcginnis@hsc.wvu.edu
rriffle@hsc.wvu.edu
mcgrewAProxyWVUH@WVUHSC.onmicrosoft.com
mmcgushin@hsc.wvu.edu
Bruce.McHam@hsc.wvu.edu
scot.mcintosh@hsc.wvu.edu
dmcintyre@hsc.wvu.edu
bmcjunkin@hsc.wvu.edu
jmcjunkin@hsc.wvu.edu
tmckeever@hsc.wvu.edu
smckendall@hsc.wvu.edu
susan.mckenrick@hsc.wvu.edu
CAMCKINLEY@hsc.wvu.edu
dmclaughlin@hsc.wvu.edu
heather.mclaughlin@hsc.wvu.edu
mark.mclaughlin@hsc.wvu.edu
smclaughlin@hsc.wvu.edu
nathanael.mcleod@hsc.wvu.edu
tmcmanus@hsc.wvu.edu
amcmillan@hsc.wvu.edu
bmcmillan@hsc.wvu.edu
mcmillenproxy@hsc.wvu.edu
jmmcmillen@hsc.wvu.edu
lmcmillen@hsc.wvu.edu
mcmillenproxy0489@WVUHSC.onmicrosoft.com
brent.mcmillion@hsc.wvu.edu
dlmcmillion@hsc.wvu.edu
kmcmillion@hsc.wvu.edu
MLMCMILLION@hsc.wvu.edu
dmcneil@hsc.wvu.edu
tmcpherson@hsc.wvu.edu
jfleshman@hsc.wvu.edu
jm0081@hsc.wvu.edu
kourtnie.mcquillen@hsc.wvu.edu
MDM@hsc.wvu.edu
mdtvconference@hsc.wvu.edu
mdtv@hsc.wvu.edu
lmeades@hsc.wvu.edu
mjmeador@hsc.wvu.edu
Carmella.Meadows@hsc.wvu.edu
Deborah.Meadows@hsc.wvu.edu
gpmeares@hsc.wvu.edu
jmears@hsc.wvu.edu
rmeckstroth@hsc.wvu.edu
km0047@WVUHSC.onmicrosoft.com
MTM@hsc.wvu.edu
medadmissions@hsc.wvu.edu
MedLeave@hsc.wvu.edu
JMEEKER1@hsc.wvu.edu
imehmi@hsc.wvu.edu
meera.mehta@hsc.wvu.edu
rashi.mehta@hsc.wvu.edu
Elizabeth.Meinert@hsc.wvu.edu
nidsy.mejiaroque@hsc.wvu.edu
mmeleady@hsc.wvu.edu
amellott@hsc.wvu.edu
kmenear@hsc.wvu.edu
amerbedone@hsc.wvu.edu
mercerproxy@hsc.wvu.edu
christopher.mercer@hsc.wvu.edu
kmercer@hsc.wvu.edu
mercerproxy1613@WVUHSC.onmicrosoft.com
aamerendino@hsc.wvu.edu
mmerzouk@hsc.wvu.edu
cmessenger@hsc.wvu.edu
ammesser@hsc.wvu.edu
pmeszaros@hsc.wvu.edu
nicki.metts@hsc.wvu.edu
alicia.meyer@hsc.wvu.edu
ashley.meyer@hsc.wvu.edu
amiah@hsc.wvu.edu
ADMICHAEL@hsc.wvu.edu
bmichael@hsc.wvu.edu
tdmichael@hsc.wvu.edu
michalskik-proxy@hsc.wvu.edu
michalskik-proxy6829@WVUHSC.onmicrosoft.com
microconfroom@hsc.wvu.edu
microcirculation@hsc.wvu.edu
microsoft@hsc.wvu.edu
microsoft1@hsc.wvu.edu
microsoft2@hsc.wvu.edu
microsoft3@hsc.wvu.edu
microsoft4@hsc.wvu.edu
TSMIDKIFF@hsc.wvu.edu
jmier@hsc.wvu.edu
migrateme1@hsc.wvu.edu
mmijuskovic@hsc.wvu.edu
lmikeo@hsc.wvu.edu
beverly.milam@hsc.wvu.edu
HBRAGG@hsc.wvu.edu
MLMILAM@hsc.wvu.edu
Bruce.Milburn@hsc.wvu.edu
walk100miles@hsc.wvu.edu
acmiller2@hsc.wvu.edu
aimiller1@hsc.wvu.edu
bmmiller@hsc.wvu.edu
bmiller@hsc.wvu.edu
ccorbett@hsc.wvu.edu
CATMILLER@hsc.wvu.edu
cmmiller@hsc.wvu.edu
Daniel.Miller1@hsc.wvu.edu
dmiller@hsc.wvu.edu
jmiller@hsc.wvu.edu
jhmiller1@hsc.wvu.edu
joshua.miller1@hsc.wvu.edu
lamiller@hsc.wvu.edu
liv.miller@hsc.wvu.edu
mark.miller1@hsc.wvu.edu
mmille52@hsc.wvu.edu
mmm0037@WVUHSC.onmicrosoft.com
mmiller@hsc.wvu.edu
romiller@hsc.wvu.edu
rgmiller@hsc.wvu.edu
sfmiller1@hsc.wvu.edu
tmiller@hsc.wvu.edu
tsmiller@hsc.wvu.edu
Zachary.Miller2@hsc.wvu.edu
millerByersProxyWVUH@WVUHSC.onmicrosoft.com
ajmillerfrost@hsc.wvu.edu
SAMILLHAM@hsc.wvu.edu
MMILLIK1@hsc.wvu.edu
amy.mills@hsc.wvu.edu
jdmills@hsc.wvu.edu
sarah.milne@hsc.wvu.edu
jminardi@hsc.wvu.edu
kminardo@hsc.wvu.edu
Samantha.Minc@wvumedicine.org
eminchau@hsc.wvu.edu
alminer@hsc.wvu.edu
fminnear@hsc.wvu.edu
1195-minolta363@hsc.wvu.edu
MIRC-CONF@hsc.wvu.edu
cbmiser@hsc.wvu.edu
RAMISRA@hsc.wvu.edu
mimitchell@hsc.wvu.edu
tmitchell@hsc.wvu.edu
amittal@hsc.wvu.edu
anne.mix@hsc.wvu.edu
Alan.Mizener@hsc.wvu.edu
mlkadmin@hsc.wvu.edu
moatsDProxyWVUH@WVUHSC.onmicrosoft.com
rmobley@hsc.wvu.edu
kmock2@hsc.wvu.edu
FRMOCNIAK@hsc.wvu.edu
rmocniak@hsc.wvu.edu
SMODI@hsc.wvu.edu
MODIFYCED@hsc.wvu.edu
kmoffett@hsc.wvu.edu
nmogge@hsc.wvu.edu
hesham.mohamed@hsc.wvu.edu
JSMOHAMED@hsc.wvu.edu
petaiah.mohan@hsc.wvu.edu
naser.moiduddin@hsc.wvu.edu
alicia.moise@hsc.wvu.edu
kmolchanoff@hsc.wvu.edu
dmolisee@hsc.wvu.edu
mamonahan@hsc.wvu.edu
dmonday@hsc.wvu.edu
amonseau@hsc.wvu.edu
MDMONTAGUE@hsc.wvu.edu
PAMONTAGUE@hsc.wvu.edu
lisa.monteville@hsc.wvu.edu
cmontgo2@hsc.wvu.edu
lmontgomery@hsc.wvu.edu
comontgomery@hsc.wvu.edu
emontgomery@hsc.wvu.edu
gm0041@hsc.wvu.edu
areynol2@hsc.wvu.edu
ahmoore@hsc.wvu.edu
camoore@hsc.wvu.edu
cemoore@hsc.wvu.edu
fletcher.moore@hsc.wvu.edu
imoore3@hsc.wvu.edu
Jennifer.Moore@hsc.wvu.edu
kathleen.moore@hsc.wvu.edu
kmoore13@hsc.wvu.edu
lmoore@hsc.wvu.edu
melissa.moore1@hsc.wvu.edu
mooremis@hsc.wvu.edu
nmdavis@hsc.wvu.edu
vamoore@hsc.wvu.edu
VNMOORE@hsc.wvu.edu
wmoore10@hsc.wvu.edu
bdmoorehead@hsc.wvu.edu
jmoorehead@hsc.wvu.edu
mooresProxyWVUH@WVUHSC.onmicrosoft.com
anvaught@hsc.wvu.edu
aeleinweber@hsc.wvu.edu
rlmoran@hsc.wvu.edu
tanya.moran@hsc.wvu.edu
wreger1@hsc.wvu.edu
moreabout@hsc.wvu.edu
jamoreland@hsc.wvu.edu
mmorela1@hsc.wvu.edu
jmorency@hsc.wvu.edu
emorgan4@hsc.wvu.edu
jlmorgan@hsc.wvu.edu
smorgan@hsc.wvu.edu
tmorise@hsc.wvu.edu
cmorley1@hsc.wvu.edu
HHICKMAN@hsc.wvu.edu
amorley@hsc.wvu.edu
ammorris1@hsc.wvu.edu
smorris@hsc.wvu.edu
tomorris@hsc.wvu.edu
LLMORRISON@hsc.wvu.edu
mary.morrison2@hsc.wvu.edu
cmortonmcswain@hsc.wvu.edu
bdmoser@hsc.wvu.edu
amoss@hsc.wvu.edu
pmoss@hsc.wvu.edu
cmott@hsc.wvu.edu
MICHELEMOUNT@hsc.wvu.edu
john.mourany@hsc.wvu.edu
amousa@hsc.wvu.edu
ymousattat@hsc.wvu.edu
Jaelyn.Mozie@hsc.wvu.edu
mph-pbe@hsc.wvu.edu
msproxy@WVUHSC.onmicrosoft.com
msstudy@hsc.wvu.edu
mthoma36proxy@hsc.wvu.edu
AMUELLE2@hsc.wvu.edu
hassan.mujahid@hsc.wvu.edu
RAMULINTI@hsc.wvu.edu
kevin.mullen@hsc.wvu.edu
kmullens@hsc.wvu.edu
cmullett@hsc.wvu.edu
mmullett@hsc.wvu.edu
rmullin2@hsc.wvu.edu
krmullins@hsc.wvu.edu
lmullin5@hsc.wvu.edu
suzanne.mundy@hsc.wvu.edu
muhamad.munir@hsc.wvu.edu
takashi.murashita@wvumedicine.org
amie.muraski@hsc.wvu.edu
carla.murgia@hsc.wvu.edu
almurphy@hsc.wvu.edu
dsmurphy@hsc.wvu.edu
tmurphy@hsc.wvu.edu
wlmurphy@hsc.wvu.edu
lmurray@hsc.wvu.edu
amurray8@hsc.wvu.edu
dmurray@hsc.wvu.edu
gmurray@hsc.wvu.edu
jessica.murray@hsc.wvu.edu
kmurray@hsc.wvu.edu
mcmurray@hsc.wvu.edu
pmurray@hsc.wvu.edu
remurray@hsc.wvu.edu
murraycProxyWVUH@WVUHSC.onmicrosoft.com
murrayJProxyWVUH@WVUHSC.onmicrosoft.com
arthur.muse@hsc.wvu.edu
kelsey.musgrove@hsc.wvu.edu
musictherapy@hsc.wvu.edu
sjmustafa@hsc.wvu.edu
hiren.muzumdar@hsc.wvu.edu
akmyers@hsc.wvu.edu
allen.myers@hsc.wvu.edu
amyers@hsc.wvu.edu
amyers14@hsc.wvu.edu
cmyers@hsc.wvu.edu
DJMYERS@hsc.wvu.edu
elmyers@hsc.wvu.edu
samuel.myers@hsc.wvu.edu
minagib@hsc.wvu.edu
savita.naik@hsc.wvu.edu
jnaim@hsc.wvu.edu
sanaime@hsc.wvu.edu
rajesh.nair@hsc.wvu.edu
dvnajar@hsc.wvu.edu
sidra.najeeb@hsc.wvu.edu
unajib@hsc.wvu.edu
Rasha.Nakity@hsc.wvu.edu
TUNANAVATI@hsc.wvu.edu
gaurav.nanda@hsc.wvu.edu
nnanda1@hsc.wvu.edu
ananjundappa@hsc.wvu.edu
syeda.naqvi@hsc.wvu.edu
karthikeyan.narayanan@hsc.wvu.edu
bnardella@hsc.wvu.edu
gnarsavage@hsc.wvu.edu
JKNARUMANCHI@hsc.wvu.edu
tnarumanchi@hsc.wvu.edu
danash@hsc.wvu.edu
jynasr@hsc.wvu.edu
layla.nasr@hsc.wvu.edu
bnass@hsc.wvu.edu
jdnasser@hsc.wvu.edu
Krupa.Nataraj@hsc.wvu.edu
anathaniel@hsc.wvu.edu
jwn0003@hsc.wvu.edu
osvaldo.navia@hsc.wvu.edu
NANAWAR@hsc.wvu.edu
carol.nay@hsc.wvu.edu
mnayeem@hsc.wvu.edu
ksnayper@hsc.wvu.edu
rnaz@hsc.wvu.edu
hanazha@hsc.wvu.edu
NBA_Conference_Room@hsc.wvu.edu
NBA_Lab_Gross_4004@hsc.wvu.edu
NBA_Lab_Gross_4006@hsc.wvu.edu
NBA_Lab_Histology@hsc.wvu.edu
NBA_Lab_SBLC@hsc.wvu.edu
obinna.ndubuizu@hsc.wvu.edu
oin0001@WVUHSC.onmicrosoft.com
shneal@hsc.wvu.edu
wneal@hsc.wvu.edu
enease@hsc.wvu.edu
lneathery@hsc.wvu.edu
kneece@hsc.wvu.edu
jason.neel@hsc.wvu.edu
gneely@hsc.wvu.edu
neelyj@hsc.wvu.edu
neeseMProxyWVUH@WVUHSC.onmicrosoft.com
isabela.negrin@hsc.wvu.edu
jneidhar@hsc.wvu.edu
lnelson@hsc.wvu.edu
thnelson@hsc.wvu.edu
sneptune@hsc.wvu.edu
lnesmith@hsc.wvu.edu
jnesselrodt@hsc.wvu.edu
knesselrodt@hsc.wvu.edu
Sydney.Nestor@hsc.wvu.edu
sarita.neupane@hsc.wvu.edu
NeuroConfRm@hsc.wvu.edu
NeurologyConferenceRoom@hsc.wvu.edu
maxwell.newby@hsc.wvu.edu
kmnewcomb@hsc.wvu.edu
snewfield@hsc.wvu.edu
atorbich@hsc.wvu.edu
cpawlak@hsc.wvu.edu
mark.newhouse@hsc.wvu.edu
jgnewman@hsc.wvu.edu
teddy.neyman@hsc.wvu.edu
pngan@hsc.wvu.edu
eynguyen@WVUHSC.onmicrosoft.com
nguyenj@hsc.wvu.edu
julian.nguyen@hsc.wvu.edu
phillip.nguyen@hsc.wvu.edu
uhnguyen@WVUHSC.onmicrosoft.com
Faraze.Niazi@hsc.wvu.edu
lnicholas@hsc.wvu.edu
matthew.nicholls@hsc.wvu.edu
ANICHOLS@hsc.wvu.edu
rnichols@hsc.wvu.edu
nnicholson@hsc.wvu.edu
pnicholson@hsc.wvu.edu
msnickasch@hsc.wvu.edu
anicola@hsc.wvu.edu
anicoloudakis@hsc.wvu.edu
honicolwala@hsc.wvu.edu
NICUreunion@hsc.wvu.edu
sniederriter@hsc.wvu.edu
lnield@hsc.wvu.edu